library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;
USE ieee.numeric_std.ALL;
entity bf6_m is
generic(Bi : integer := 16);
Port (     por   : in std_logic;
	        a2_r  : in std_logic_vector(Bi - 1 downto 0);
	        a2_i  : in std_logic_vector(Bi - 1 downto 0);
           a21_r : in std_logic_vector(Bi - 1 downto 0);
	        a21_i : in std_logic_vector(Bi - 1 downto 0);
			  i     : in std_logic;
			  i1    : in std_logic;
			  i4    : in std_logic;
			  b2_r  : out std_logic_vector(Bi-1 downto 0);
			  b2_i  : out std_logic_vector(Bi-1 downto 0);
			  b21_r : out std_logic_vector(Bi-1 downto 0);
			  b21_i : out std_logic_vector(Bi-1 downto 0)
			 );
end bf6_m;
architecture Behavioral of bf6_m is
begin
process(por,i4)
begin
  if(por='1') then
      b2_r <=   (others => '0'); 
		b2_i <=   (others => '0'); 
		b21_r <=  (others => '0'); 
		b21_i <=  (others => '0'); 

  elsif(i4 = '1') then
		if i = '0'  then
			b2_r  <= (a2_r) ;
			b2_i  <= (a2_i) ;
			b21_r <= (a21_r) ;
			b21_i <= (a21_i) ;
		else
			if i1 = '1'  then
				b2_r <=  (a21_r) - (a2_r) ;
				b2_i <=  (a21_i) - (a2_i) ;
				b21_r <= (a21_r) + (a2_r);
				b21_i <= (a21_i) + (a2_i);
			else
				b2_r  <= (a21_r)  - (a2_i) ; 
				b2_i  <= (a21_i)  + (a2_r) ; 
				b21_r <= (a21_r)  + (a2_i); 
				b21_i <= (a21_i)  - (a2_r) ; 
			end if;
		end if;
   end if;
end process;
end Behavioral;